module axi_memory();
endmodule
